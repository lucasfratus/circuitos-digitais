CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 1 90 10
163 80 1598 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
331 176 444 273
9437202 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 24 90 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 CLK
-10 -31 11 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6986 0 0
2
45360.7 0
0
13 Logic Switch~
5 80 93 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 PR
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8745 0 0
2
45360.7 1
0
9 2-In AND~
219 585 782 0 3 22
0 5 3 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9592 0 0
2
45360.7 2
0
9 2-In AND~
219 439 746 0 3 22
0 3 6 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8748 0 0
2
45360.7 3
0
6 74112~
219 672 712 0 7 32
0 10 7 11 3 4 6 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U6A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 6 0
1 U
7168 0 0
2
45360.7 4
0
6 74112~
219 513 686 0 7 32
0 10 8 11 3 4 19 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U5B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 5 0
1 U
631 0 0
2
45360.7 5
0
6 74112~
219 349 664 0 7 32
0 10 10 11 4 4 20 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U5A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 5 0
1 U
9466 0 0
2
45360.7 6
0
12 Hex Display~
7 938 117 0 18 19
10 3 5 9 21 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3266 0 0
2
45360.7 7
0
12 Hex Display~
7 1003 117 0 18 19
10 2 12 13 11 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7693 0 0
2
45360.7 8
0
5 7415~
219 718 509 0 4 22
0 13 12 2 17
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 4 0
1 U
3723 0 0
2
45360.7 9
0
9 2-In AND~
219 516 491 0 3 22
0 12 2 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3440 0 0
2
45360.7 10
0
9 2-In AND~
219 320 454 0 3 22
0 2 14 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6263 0 0
2
45360.7 11
0
7 Pulser~
4 65 336 0 10 12
0 22 23 18 24 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4900 0 0
2
45360.7 12
0
6 74112~
219 792 273 0 7 32
0 10 17 18 2 4 14 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 2 0
1 U
8783 0 0
2
45360.7 13
0
6 74112~
219 652 273 0 7 32
0 10 15 18 15 4 25 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3221 0 0
2
45360.7 14
0
6 74112~
219 502 272 0 7 32
0 10 16 18 2 4 26 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3215 0 0
2
45360.7 15
0
6 74112~
219 348 265 0 7 32
0 10 10 18 18 4 2 2
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
7903 0 0
2
45360.7 16
0
54
4 0 2 0 0 8192 0 14 0 0 25 3
768 255
762 255
762 190
2 0 3 0 0 8192 0 3 0 0 3 3
561 791
532 791
532 703
4 0 3 0 0 12288 0 5 0 0 11 5
648 694
552 694
552 703
425 703
425 668
4 0 4 0 0 8192 0 7 0 0 7 3
325 646
294 646
294 728
5 0 4 0 0 0 0 6 0 0 7 2
513 698
513 728
5 0 4 0 0 0 0 7 0 0 7 2
349 676
349 728
5 0 4 0 0 8192 0 5 0 0 38 4
672 724
672 728
184 728
184 401
1 0 5 0 0 8192 0 3 0 0 14 3
561 773
549 773
549 650
2 6 6 0 0 12416 0 4 5 0 0 6
415 755
406 755
406 765
710 765
710 694
702 694
3 2 7 0 0 8320 0 3 5 0 0 4
606 782
634 782
634 676
648 676
4 0 3 0 0 0 0 6 0 0 16 2
489 668
387 668
3 2 8 0 0 8320 0 4 6 0 0 4
460 746
475 746
475 650
489 650
7 3 9 0 0 8320 0 5 8 0 0 3
696 676
935 676
935 141
7 2 5 0 0 8320 0 6 8 0 0 3
537 650
941 650
941 141
0 1 3 0 0 4224 0 0 8 16 0 3
387 628
947 628
947 141
1 7 3 0 0 0 0 4 7 0 0 4
415 737
387 737
387 628
373 628
2 0 10 0 0 8192 0 7 0 0 23 3
325 628
311 628
311 595
3 0 11 0 0 8192 0 5 0 0 20 3
642 685
621 685
621 578
3 0 11 0 0 0 0 6 0 0 20 3
483 659
471 659
471 578
3 0 11 0 0 12416 0 7 0 0 28 5
319 637
291 637
291 578
881 578
881 237
1 0 10 0 0 0 0 7 0 0 23 2
349 601
349 595
1 0 10 0 0 0 0 6 0 0 23 2
513 623
513 595
0 1 10 0 0 8192 0 0 5 54 0 4
108 139
108 595
672 595
672 649
4 0 2 0 0 4096 0 16 0 0 25 3
478 254
390 254
390 229
0 1 2 0 0 12416 0 0 9 33 0 5
377 229
392 229
392 190
1012 190
1012 141
0 2 12 0 0 12416 0 0 9 40 0 5
542 236
555 236
555 205
1006 205
1006 141
0 3 13 0 0 12416 0 0 9 30 0 5
710 237
712 237
712 216
1000 216
1000 141
7 4 11 0 0 0 0 14 9 0 0 3
816 237
994 237
994 141
1 0 2 0 0 0 0 12 0 0 33 3
296 445
296 416
377 416
1 7 13 0 0 0 0 10 15 0 0 6
694 500
688 500
688 289
710 289
710 237
676 237
2 0 2 0 0 0 0 11 0 0 33 2
492 500
377 500
6 0 2 0 0 0 0 17 0 0 33 2
378 247
377 247
3 7 2 0 0 0 0 10 17 0 0 4
694 518
377 518
377 229
372 229
2 6 14 0 0 12416 0 12 14 0 0 6
296 463
275 463
275 370
830 370
830 255
822 255
5 0 4 0 0 0 0 15 0 0 38 2
652 285
652 401
5 0 4 0 0 0 0 16 0 0 38 2
502 284
502 401
5 0 4 0 0 0 0 17 0 0 38 2
348 277
348 401
1 5 4 0 0 8320 0 1 14 0 0 4
24 102
24 401
792 401
792 285
1 0 12 0 0 0 0 11 0 0 40 3
492 482
492 437
542 437
2 7 12 0 0 0 0 10 16 0 0 4
694 509
542 509
542 236
526 236
4 0 15 0 0 4096 0 15 0 0 42 2
628 255
618 255
3 2 15 0 0 8320 0 11 15 0 0 4
537 491
618 491
618 237
628 237
2 3 16 0 0 8320 0 16 12 0 0 4
478 236
407 236
407 454
341 454
4 2 17 0 0 8320 0 10 14 0 0 4
739 509
748 509
748 237
768 237
4 0 18 0 0 8192 0 17 0 0 49 3
324 247
262 247
262 327
3 0 18 0 0 8192 0 17 0 0 49 3
318 238
295 238
295 327
3 0 18 0 0 0 0 16 0 0 49 3
472 245
438 245
438 327
3 0 18 0 0 0 0 15 0 0 49 3
622 246
597 246
597 327
3 3 18 0 0 4224 0 13 14 0 0 4
89 327
754 327
754 246
762 246
2 0 10 0 0 0 0 17 0 0 54 3
324 229
308 229
308 137
1 0 10 0 0 0 0 17 0 0 54 2
348 202
348 137
1 0 10 0 0 0 0 16 0 0 54 2
502 209
502 137
1 0 10 0 0 0 0 15 0 0 54 2
652 210
652 137
1 1 10 0 0 8320 0 14 2 0 0 4
792 210
792 137
80 137
80 105
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
