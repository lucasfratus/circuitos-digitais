CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 910 30 80 10
81 80 1598 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
249 176 362 273
42991634 0
0
6 Title:
5 Name:
0
0
0
66
13 Logic Switch~
5 19 1319 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 OE
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90115e-315 0
0
13 Logic Switch~
5 21 1236 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 RD
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90115e-315 0
0
13 Logic Switch~
5 20 1166 0 1 11
0 21
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 CS
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.90115e-315 0
0
13 Logic Switch~
5 22 35 0 1 11
0 6
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.90115e-315 0
0
13 Logic Switch~
5 81 33 0 1 11
0 8
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 A0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90115e-315 0
0
13 Logic Switch~
5 1156 104 0 1 11
0 11
0
0 0 21344 180
2 0V
-7 -16 7 -8
2 I1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.90115e-315 0
0
13 Logic Switch~
5 1153 147 0 1 11
0 44
0
0 0 21344 180
2 0V
-7 -16 7 -8
2 I0
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.90115e-315 0
0
13 Logic Switch~
5 1160 60 0 1 11
0 52
0
0 0 21344 180
2 0V
-7 -16 7 -8
2 I2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 166 706 0 3 22
0 7 6 5
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U23A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
4747 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 167 506 0 3 22
0 8 9 4
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U20D
-18 -26 10 -18
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
972 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 164 955 0 3 22
0 8 6 3
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U20C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
3472 0 0
2
5.90115e-315 0
0
9 Inverter~
13 106 99 0 2 22
0 8 7
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 U14F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
9998 0 0
2
5.90115e-315 0
0
9 Inverter~
13 47 102 0 2 22
0 6 9
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 U14E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
3536 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 170 308 0 3 22
0 7 9 10
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U20B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
4597 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 1008 1373 0 1 2
10 12
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 D0
14 0 28 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 694 1378 0 1 2
10 13
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 D1
14 0 28 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 411 1370 0 1 2
10 14
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 D2
14 0 28 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90115e-315 0
0
10 Buffer 3S~
219 695 1298 0 3 22
0 15 17 13
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U22C
14 -5 42 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
9323 0 0
2
5.90115e-315 0
0
10 Buffer 3S~
219 1009 1295 0 3 22
0 18 17 12
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U22B
14 -5 42 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
317 0 0
2
5.90115e-315 0
0
10 Buffer 3S~
219 412 1291 0 3 22
0 16 17 14
0
0 0 608 270
8 BUFFER3S
-27 -51 29 -43
4 U22A
14 -5 42 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3108 0 0
2
5.90115e-315 0
0
5 7415~
219 247 1309 0 4 22
0 20 21 19 17
0
0 0 608 0
6 74LS15
-21 -28 21 -20
4 U21A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 9 0
1 U
4299 0 0
2
5.90115e-315 0
0
9 Inverter~
13 199 1136 0 2 22
0 20 22
0
0 0 608 90
6 74LS04
-21 -19 21 -11
4 U14C
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
9672 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 194 1058 0 3 22
0 21 22 2
0
0 0 608 90
6 74LS08
-21 -24 21 -16
4 U20A
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
7876 0 0
2
5.90115e-315 0
0
8 4-In OR~
219 1004 1131 0 5 22
0 23 24 25 26 18
0
0 0 608 270
4 4072
-14 -24 14 -16
4 U19A
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
6369 0 0
2
5.90115e-315 0
0
8 4-In OR~
219 689 1133 0 5 22
0 27 28 29 30 15
0
0 0 608 270
4 4072
-14 -24 14 -16
4 U18B
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
9172 0 0
2
5.90115e-315 0
0
8 4-In OR~
219 408 1130 0 5 22
0 31 32 33 34 16
0
0 0 608 270
4 4072
-14 -24 14 -16
4 U18A
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
7100 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 949 862 0 1 2
10 37
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 647 858 0 1 2
10 38
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 987 995 0 3 22
0 37 3 26
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U17D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
961 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 655 978 0 3 22
0 38 3 30
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U17C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3178 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 380 976 0 3 22
0 39 3 34
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U17B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3409 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 230 920 0 3 22
0 2 3 35
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U17A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3951 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 948 622 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 680 745 0 3 22
0 41 5 29
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U16D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3780 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 397 739 0 3 22
0 42 5 33
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U16C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9265 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 1002 747 0 3 22
0 40 5 25
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U16B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9442 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 231 669 0 3 22
0 2 5 36
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9424 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 238 460 0 3 22
0 2 4 43
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U15D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9968 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 941 397 0 1 2
10 45
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 1019 542 0 3 22
0 45 4 24
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U15C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8464 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 642 613 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 702 533 0 3 22
0 46 4 28
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U15B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3171 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 664 399 0 1 2
10 46
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 424 534 0 3 22
0 47 4 32
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U15A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6435 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 664 181 0 1 2
10 48
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 733 350 0 3 22
0 48 10 27
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U13D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
6874 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 964 180 0 1 2
10 51
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 1034 356 0 3 22
0 51 10 23
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U13C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
34 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 240 254 0 3 22
0 2 10 49
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
969 0 0
2
5.90115e-315 0
0
9 2-In AND~
219 452 350 0 3 22
0 50 10 31
0
0 0 608 270
6 74LS08
-21 -24 21 -16
4 U13A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8402 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 374 858 0 1 2
10 39
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 373 185 0 1 2
10 50
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 373 401 0 1 2
10 47
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
5.90115e-315 0
0
14 Logic Display~
6 372 615 0 1 2
10 42
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 845 916 0 4 9
0 44 35 53 37
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U12
-10 -55 11 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6357 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 575 912 0 4 9
0 11 35 54 38
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U11
-10 -55 11 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
319 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 306 914 0 4 9
0 52 35 55 39
0
0 0 4704 0
3 DFF
-10 -53 11 -45
3 U10
-10 -55 11 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3976 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 862 676 0 4 9
0 44 36 56 40
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U9
-7 -56 7 -48
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7634 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 585 669 0 4 9
0 11 36 57 41
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U8
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
523 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 321 668 0 4 9
0 52 36 58 42
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U7
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6748 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 864 452 0 4 9
0 44 43 59 45
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6901 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 588 455 0 4 9
0 11 43 60 46
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U5
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
842 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 318 453 0 4 9
0 52 43 61 47
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U4
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3277 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 856 233 0 4 9
0 44 49 62 51
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4212 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 600 235 0 4 9
0 11 49 63 48
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4720 0 0
2
5.90115e-315 0
0
12 D Flip-Flop~
219 316 237 0 4 9
0 52 49 64 50
0
0 0 4704 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5551 0 0
2
5.90115e-315 0
0
105
1 0 2 0 0 4096 0 37 0 0 43 2
207 660
193 660
2 0 3 0 0 8192 0 32 0 0 7 3
206 929
200 929
200 955
0 2 4 0 0 4096 0 0 38 16 0 3
206 506
206 469
214 469
0 2 5 0 0 4096 0 0 37 10 0 3
202 706
202 678
207 678
2 0 3 0 0 0 0 31 0 0 7 2
369 954
369 955
2 0 3 0 0 0 0 30 0 0 7 2
644 956
644 955
3 2 3 0 0 4224 0 11 29 0 0 3
185 955
976 955
976 973
2 0 5 0 0 0 0 34 0 0 10 2
669 723
669 706
2 0 5 0 0 0 0 35 0 0 10 2
386 717
386 706
3 2 5 0 0 4224 0 9 36 0 0 3
187 706
991 706
991 725
2 0 6 0 0 4096 0 9 0 0 25 2
142 715
23 715
1 0 2 0 0 0 0 32 0 0 43 2
206 911
193 911
1 0 7 0 0 8320 0 9 0 0 21 3
142 697
109 697
109 299
2 0 4 0 0 0 0 42 0 0 16 2
691 511
691 506
2 0 4 0 0 0 0 44 0 0 16 3
413 512
413 506
411 506
2 3 4 0 0 8320 0 40 10 0 0 3
1008 520
1008 506
188 506
0 1 8 0 0 4096 0 0 10 23 0 2
81 497
143 497
0 2 9 0 0 4224 0 0 10 20 0 3
50 315
50 515
143 515
1 0 2 0 0 8192 0 49 0 0 43 4
216 245
192 245
192 451
193 451
2 2 9 0 0 0 0 13 14 0 0 3
50 120
50 317
146 317
2 1 7 0 0 0 0 12 14 0 0 3
109 117
109 299
146 299
1 0 8 0 0 0 0 12 0 0 23 3
109 81
109 59
81 59
1 1 8 0 0 8320 0 11 5 0 0 3
140 946
81 946
81 45
1 0 6 0 0 0 0 13 0 0 25 3
50 84
50 59
22 59
1 2 6 0 0 4224 0 4 11 0 0 5
22 47
22 679
23 679
23 964
140 964
3 2 10 0 0 12416 0 14 48 0 0 5
191 308
217 308
217 307
1023 307
1023 334
1 1 11 0 0 8320 0 6 56 0 0 4
1142 104
508 104
508 876
551 876
1 3 12 0 0 4224 0 15 19 0 0 2
1008 1359
1008 1311
1 3 13 0 0 4224 0 16 18 0 0 2
694 1364
694 1314
1 3 14 0 0 4224 0 17 20 0 0 2
411 1356
411 1307
1 5 15 0 0 4224 0 18 25 0 0 4
694 1284
694 1166
692 1166
692 1163
1 5 16 0 0 4224 0 20 26 0 0 2
411 1277
411 1160
2 0 17 0 0 8192 0 20 0 0 36 3
400 1292
366 1292
366 1240
2 0 17 0 0 8192 0 18 0 0 36 3
683 1299
657 1299
657 1240
1 5 18 0 0 4224 0 19 24 0 0 4
1008 1281
1008 1176
1007 1176
1007 1161
2 4 17 0 0 12416 0 19 21 0 0 6
997 1296
962 1296
962 1240
276 1240
276 1309
268 1309
3 1 19 0 0 4224 0 21 1 0 0 4
223 1318
40 1318
40 1319
31 1319
1 0 20 0 0 4096 0 2 0 0 40 2
33 1236
115 1236
2 0 21 0 0 4096 0 21 0 0 41 3
223 1309
75 1309
75 1166
1 1 20 0 0 4224 0 21 22 0 0 5
223 1300
115 1300
115 1236
202 1236
202 1154
1 1 21 0 0 8320 0 23 3 0 0 3
184 1079
184 1166
32 1166
2 2 22 0 0 4224 0 22 23 0 0 2
202 1118
202 1079
3 1 2 0 0 4224 0 23 38 0 0 3
193 1034
193 451
214 451
1 3 23 0 0 4224 0 24 48 0 0 7
1020 1111
1020 800
1036 800
1036 563
1038 563
1038 379
1032 379
2 3 24 0 0 4224 0 24 40 0 0 6
1011 1111
1011 790
1020 790
1020 567
1017 567
1017 565
3 3 25 0 0 12416 0 24 36 0 0 6
1002 1111
1002 1033
1006 1033
1006 794
1000 794
1000 770
4 3 26 0 0 4224 0 24 29 0 0 4
993 1111
993 1037
985 1037
985 1018
1 3 27 0 0 12416 0 25 46 0 0 7
705 1113
705 1039
712 1039
712 571
732 571
732 373
731 373
2 3 28 0 0 12416 0 25 42 0 0 4
696 1113
696 1031
700 1031
700 556
3 3 29 0 0 12416 0 25 34 0 0 4
687 1113
687 1026
678 1026
678 768
4 3 30 0 0 4224 0 25 30 0 0 4
678 1113
678 1030
653 1030
653 1001
2 0 10 0 0 0 0 50 0 0 26 2
441 328
441 307
2 0 10 0 0 0 0 46 0 0 26 2
722 328
722 307
1 3 31 0 0 12416 0 26 50 0 0 4
424 1110
424 1070
450 1070
450 373
2 3 32 0 0 12416 0 26 44 0 0 6
415 1110
415 1057
423 1057
423 565
422 565
422 557
3 3 33 0 0 4224 0 26 35 0 0 4
406 1110
406 790
395 790
395 762
4 3 34 0 0 12416 0 26 31 0 0 4
397 1110
397 1072
378 1072
378 999
2 0 35 0 0 8192 0 56 0 0 62 3
551 894
539 894
539 921
2 0 36 0 0 4096 0 59 0 0 73 3
561 651
542 651
542 669
2 0 36 0 0 0 0 60 0 0 73 3
297 650
289 650
289 669
2 0 35 0 0 0 0 57 0 0 62 3
282 896
255 896
255 921
3 2 35 0 0 12416 0 32 55 0 0 6
251 920
255 920
255 921
813 921
813 898
821 898
1 0 37 0 0 0 0 27 0 0 65 2
949 880
949 880
1 0 38 0 0 0 0 28 0 0 66 2
647 876
647 876
1 4 37 0 0 8320 0 29 55 0 0 3
994 973
994 880
869 880
1 4 38 0 0 4224 0 30 56 0 0 3
662 956
662 876
599 876
1 1 39 0 0 4224 0 31 51 0 0 4
387 954
387 878
374 878
374 876
1 0 40 0 0 0 0 33 0 0 69 2
948 640
948 640
1 4 40 0 0 8320 0 36 58 0 0 3
1009 725
1009 640
886 640
1 0 41 0 0 4096 0 41 0 0 71 2
642 631
642 633
1 4 41 0 0 4224 0 34 59 0 0 3
687 723
687 633
609 633
1 1 42 0 0 4224 0 35 54 0 0 3
404 717
404 633
372 633
3 2 36 0 0 4224 0 37 58 0 0 4
252 669
830 669
830 658
838 658
2 0 43 0 0 8192 0 62 0 0 76 3
564 437
546 437
546 460
0 2 43 0 0 4096 0 0 63 76 0 3
284 460
284 435
294 435
3 2 43 0 0 4224 0 38 61 0 0 4
259 460
832 460
832 434
840 434
1 0 44 0 0 8192 0 58 0 0 102 3
838 640
838 637
777 637
1 0 45 0 0 4096 0 39 0 0 79 2
941 415
941 416
1 4 45 0 0 8320 0 40 61 0 0 3
1026 520
1026 416
888 416
0 2 10 0 0 0 0 0 49 26 0 3
212 307
212 263
216 263
1 0 46 0 0 8192 0 43 0 0 82 3
664 417
663 417
663 420
1 4 46 0 0 4224 0 42 62 0 0 5
709 511
709 420
663 420
663 419
612 419
1 0 44 0 0 4096 0 61 0 0 102 2
840 416
777 416
1 1 47 0 0 4224 0 44 53 0 0 3
431 512
431 419
373 419
1 0 48 0 0 0 0 45 0 0 86 2
664 199
664 199
4 1 48 0 0 8320 0 65 46 0 0 3
624 199
740 199
740 328
2 0 49 0 0 8192 0 65 0 0 92 3
576 217
561 217
561 254
2 0 49 0 0 0 0 66 0 0 92 3
292 219
286 219
286 254
1 1 50 0 0 4224 0 50 52 0 0 4
459 328
459 201
373 201
373 203
1 0 51 0 0 8192 0 47 0 0 91 3
964 198
964 197
988 197
1 4 51 0 0 8320 0 48 64 0 0 3
1041 334
1041 197
880 197
3 2 49 0 0 4224 0 49 64 0 0 4
261 254
824 254
824 215
832 215
1 0 44 0 0 0 0 64 0 0 102 2
832 197
777 197
4 1 39 0 0 0 0 57 51 0 0 3
330 878
374 878
374 876
1 4 42 0 0 0 0 54 60 0 0 4
372 633
359 633
359 632
345 632
4 1 47 0 0 0 0 63 53 0 0 3
342 417
373 417
373 419
4 1 50 0 0 0 0 66 52 0 0 3
340 201
373 201
373 203
1 0 52 0 0 4096 0 66 0 0 101 2
292 201
260 201
1 0 52 0 0 0 0 63 0 0 101 4
294 417
275 417
275 418
260 418
1 0 52 0 0 0 0 60 0 0 101 4
297 632
275 632
275 633
259 633
1 1 52 0 0 12416 0 57 8 0 0 5
282 878
259 878
259 63
1146 63
1146 60
1 1 44 0 0 8320 0 55 7 0 0 4
821 880
777 880
777 147
1139 147
1 0 11 0 0 0 0 65 0 0 27 2
576 199
508 199
1 0 11 0 0 0 0 62 0 0 27 2
564 419
508 419
1 0 11 0 0 0 0 59 0 0 27 4
561 633
523 633
523 632
508 632
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
